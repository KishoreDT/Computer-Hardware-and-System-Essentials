* C:\POE\EX3.sch

* Schematics Version 9.1 - Web Update 1
* Mon May 16 13:50:58 2022



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "EX3.net"
.INC "EX3.als"


.probe


.END
