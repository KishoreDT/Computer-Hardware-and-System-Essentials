* C:\POE\EX5.sch

* Schematics Version 9.1 - Web Update 1
* Mon May 16 21:07:28 2022



** Analysis setup **
.tran 0ns 5ms
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "EX5.net"
.INC "EX5.als"


.probe


.END
