* C:\POE\EX4.sch

* Schematics Version 9.1 - Web Update 1
* Mon May 16 13:57:51 2022



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "EX4.net"
.INC "EX4.als"


.probe


.END
